//------------------------------------------------------//
//- Advanced Digital IC Design                          //
//-                                                     //
//- Exercise: Design a FSK Modem                        //
//------------------------------------------------------//
`timescale 1ns/1ps
`include "MONITOR.v"
`include "PFD.v"
`include "CONTROLLER.v"
`include "dco_model.v"
`include "frequency_div.v"
module TOP;
wire [131 : 0] DCO_CODE;
wire [2 : 0] M;
MONITOR    MONITOR(.reset(RESET),
                   .reset_(RESET_),
                   .ref_clk(REF_CLK),
                   .m(M)
                   );
PFD        PFD(.ref_clk(REF_CLK),
               .fb(Out_divM),
               .flagu(FLAGU),
               .flagd(FLAGD)
               );
CONTROLLER CONTROLLER(.reset(RESET),
                      .p_up(FLAGU),
                      .p_down(FLAGD), 
                      .dco_code(DCO_CODE),
                      .freq_lock(FREQ_LOCK),
                      .polarity(POLARITY)
                      );
dco_model  dco_model(.reset_(RESET_),   
                  .en_0(DCO_CODE[0]),
                  .en_1(DCO_CODE[1]), 
                  .en_2(DCO_CODE[2]), 
                  .en_3(DCO_CODE[3]),
                  .en_4(DCO_CODE[4]),
                  .en_5(DCO_CODE[5]), 
                  .en_6(DCO_CODE[6]), 
                  .en_7(DCO_CODE[7]),
                  .en_8(DCO_CODE[8]),
                  .en_9(DCO_CODE[9]), 
                  .en_10(DCO_CODE[10]), 
                  .en_11(DCO_CODE[11]),
                  .en_12(DCO_CODE[12]),
                  .en_13(DCO_CODE[13]), 
                  .en_14(DCO_CODE[14]), 
                  .en_15(DCO_CODE[15]), 
                  .en_16(DCO_CODE[16]),
                  .en_17(DCO_CODE[17]), 
                  .en_18(DCO_CODE[18]), 
                  .en_19(DCO_CODE[19]),
                  .en_20(DCO_CODE[20]),
                  .en_21(DCO_CODE[21]), 
                  .en_22(DCO_CODE[22]), 
                  .en_23(DCO_CODE[23]), 
                  .en_24(DCO_CODE[24]),
                  .en_25(DCO_CODE[25]), 
                  .en_26(DCO_CODE[26]), 
                  .en_27(DCO_CODE[27]),
                  .en_28(DCO_CODE[28]),
                  .en_29(DCO_CODE[29]), 
                  .en_30(DCO_CODE[30]), 
                  .en_31(DCO_CODE[31]), 
                  .en_32(DCO_CODE[32]),
                  .en_33(DCO_CODE[33]), 
                  .en_34(DCO_CODE[34]), 
                  .en_35(DCO_CODE[35]),
                  .en_36(DCO_CODE[36]),
                  .en_37(DCO_CODE[37]), 
                  .en_38(DCO_CODE[38]), 
                  .en_39(DCO_CODE[39]), 
                  .en_40(DCO_CODE[40]),
                  .en_41(DCO_CODE[41]), 
                  .en_42(DCO_CODE[42]), 
                  .en_43(DCO_CODE[43]),
                  .en_44(DCO_CODE[44]),
                  .en_45(DCO_CODE[45]), 
                  .en_46(DCO_CODE[46]), 
                  .en_47(DCO_CODE[47]),
                  .en_48(DCO_CODE[48]),
                  .en_49(DCO_CODE[49]), 
                  .en_50(DCO_CODE[50]), 
                  .en_51(DCO_CODE[51]),
                  .en_52(DCO_CODE[52]),
                  .en_53(DCO_CODE[53]), 
                  .en_54(DCO_CODE[54]), 
                  .en_55(DCO_CODE[55]), 
                  .en_56(DCO_CODE[56]),
                  .en_57(DCO_CODE[57]), 
                  .en_58(DCO_CODE[58]), 
                  .en_59(DCO_CODE[59]),
                  .en_60(DCO_CODE[60]),
                  .en_61(DCO_CODE[61]), 
                  .en_62(DCO_CODE[62]), 
                  .en_63(DCO_CODE[63]), 
                  .en_64(DCO_CODE[64]),
                  .en_65(DCO_CODE[65]), 
                  .en_66(DCO_CODE[66]), 
                  .en_67(DCO_CODE[67]),
                  .en_68(DCO_CODE[68]),
                  .en_69(DCO_CODE[69]), 
                  .en_70(DCO_CODE[70]), 
                  .en_71(DCO_CODE[71]), 
                  .en_72(DCO_CODE[72]),
                  .en_73(DCO_CODE[73]), 
                  .en_74(DCO_CODE[74]), 
                  .en_75(DCO_CODE[75]),
                  .en_76(DCO_CODE[76]),
                  .en_77(DCO_CODE[77]), 
                  .en_78(DCO_CODE[78]), 
                  .en_79(DCO_CODE[79]),
                  .en_80(DCO_CODE[80]),
                  .en_81(DCO_CODE[81]), 
                  .en_82(DCO_CODE[82]), 
                  .en_83(DCO_CODE[83]),
                  .en_84(DCO_CODE[84]),
                  .en_85(DCO_CODE[85]), 
                  .en_86(DCO_CODE[86]), 
                  .en_87(DCO_CODE[87]), 
                  .en_88(DCO_CODE[88]),
                  .en_89(DCO_CODE[89]), 
                  .en_90(DCO_CODE[90]), 
                  .en_91(DCO_CODE[91]),
                  .en_92(DCO_CODE[92]),
                  .en_93(DCO_CODE[93]), 
                  .en_94(DCO_CODE[94]), 
                  .en_95(DCO_CODE[95]), 
                  .en_96(DCO_CODE[96]),
                  .en_97(DCO_CODE[97]), 
                  .en_98(DCO_CODE[98]), 
                  .en_99(DCO_CODE[99]),
                  .en_100(DCO_CODE[100]),
                  .en_101(DCO_CODE[101]), 
                  .en_102(DCO_CODE[102]), 
                  .en_103(DCO_CODE[103]), 
                  .en_104(DCO_CODE[104]),
                  .en_105(DCO_CODE[105]), 
                  .en_106(DCO_CODE[106]), 
                  .en_107(DCO_CODE[107]),
                  .en_108(DCO_CODE[108]),
                  .en_109(DCO_CODE[109]), 
                  .en_110(DCO_CODE[110]), 
                  .en_111(DCO_CODE[111]), 
                  .en_112(DCO_CODE[112]),
                  .en_113(DCO_CODE[113]), 
                  .en_114(DCO_CODE[114]), 
                  .en_115(DCO_CODE[115]),
                  .en_116(DCO_CODE[116]),
                  .en_117(DCO_CODE[117]), 
                  .en_118(DCO_CODE[118]), 
                  .en_119(DCO_CODE[119]),
                  .en_120(DCO_CODE[120]),
                  .en_121(DCO_CODE[121]), 
                  .en_122(DCO_CODE[122]), 
                  .en_123(DCO_CODE[123]), 
                  .en_124(DCO_CODE[124]),
                  .en_125(DCO_CODE[125]), 
                  .en_126(DCO_CODE[126]), 
                  .en_127(DCO_CODE[127]),
                  .en_128(DCO_CODE[128]),
                  .en_129(DCO_CODE[129]),
                  .en_130(DCO_CODE[130]),
                  .en_131(DCO_CODE[131]),              
                  .dco_out(OUT_CLK)
                );
frequency_div frequency_div( .n(M),
                           .ref_clk(OUT_CLK),
                           .clk_count(CLK_COUNT),
                           .clk_divn(Out_divM),
                           .reset(RESET)
                           );

endmodule